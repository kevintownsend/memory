module rr_testbench;
initial begin
    $display("hello world");
    $finish;
end
endmodule

module rr_testbench;
// TODO: clock
//signal i;
//reg clk;
//reg [0 : 3] wr;
//wire [5 : 0] wr_addr [0 : INPUTS];

//timstamp_rr dut(clk, wr, wr_addr);

initial begin
    $display("hello world");

    $finish;
end
endmodule
